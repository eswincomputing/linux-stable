--signal declaration from Document Version 1.1.2
 signal SwRegister_sw_vcmd_hw_id : std_logic_vector(15 downto 0);
 signal SwRegister_sw_vcmd_hw_version : std_logic_vector(15 downto 0);
 signal SwRegister_sw_vcmd_hw_build_date : std_logic_vector(31 downto 0);
 signal SwRegister_sw_vcmd_ext_abn_int_src_vcd_mmu : std_logic;
 signal SwRegister_sw_vcmd_ext_abn_int_src_vcd_l2cache : std_logic;
 signal SwRegister_sw_vcmd_ext_abn_int_src_vcd_dec400 : std_logic;
 signal SwRegister_sw_vcmd_ext_abn_int_src_vcd : std_logic;
 signal SwRegister_sw_vcmd_ext_abn_int_src_cutree_mmu : std_logic;
 signal SwRegister_sw_vcmd_ext_abn_int_src_vce_mmu : std_logic;
 signal SwRegister_sw_vcmd_ext_abn_int_src_vce_l2cache : std_logic;
 signal SwRegister_sw_vcmd_ext_abn_int_src_vce_dec400 : std_logic;
 signal SwRegister_sw_vcmd_ext_abn_int_src_cutree : std_logic;
 signal SwRegister_sw_vcmd_ext_abn_int_src_vce : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_vcd_mmu : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_vcd_l2cache : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_vcd_dec400 : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_vcd : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_cutree_mmu : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_vce_mmu : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_vce_l2cache : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_vce_dec400 : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_cutree : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_vce : std_logic;
 signal SwRegister_sw_vcmd_exe_cmdbuf_count : std_logic_vector(31 downto 0);
 signal SwRegister_sw_vcmd_executing_cmd : std_logic_vector(31 downto 0);
 signal SwRegister_sw_vcmd_executing_cmd_msb : std_logic_vector(31 downto 0);
 signal SwRegister_sw_vcmd_axi_total_ar_len : std_logic_vector(31 downto 0);
 signal SwRegister_sw_vcmd_axi_total_r : std_logic_vector(31 downto 0);
 signal SwRegister_sw_vcmd_axi_total_ar : std_logic_vector(31 downto 0);
 signal SwRegister_sw_vcmd_axi_total_r_last : std_logic_vector(31 downto 0);
 signal SwRegister_sw_vcmd_axi_total_aw_len : std_logic_vector(31 downto 0);
 signal SwRegister_sw_vcmd_axi_total_w : std_logic_vector(31 downto 0);
 signal SwRegister_sw_vcmd_axi_total_aw : std_logic_vector(31 downto 0);
 signal SwRegister_sw_vcmd_axi_total_w_last : std_logic_vector(31 downto 0);
 signal SwRegister_sw_vcmd_axi_total_b : std_logic_vector(31 downto 0);
 signal SwRegister_sw_vcmd_axi_ar_valid : std_logic;
 signal SwRegister_sw_vcmd_axi_ar_ready : std_logic;
 signal SwRegister_sw_vcmd_axi_r_valid : std_logic;
 signal SwRegister_sw_vcmd_axi_r_ready : std_logic;
 signal SwRegister_sw_vcmd_axi_aw_valid : std_logic;
 signal SwRegister_sw_vcmd_axi_aw_ready : std_logic;
 signal SwRegister_sw_vcmd_axi_w_valid : std_logic;
 signal SwRegister_sw_vcmd_axi_w_ready : std_logic;
 signal SwRegister_sw_vcmd_axi_b_valid : std_logic;
 signal SwRegister_sw_vcmd_axi_b_ready : std_logic;
 signal SwRegister_sw_vcmd_work_state : std_logic_vector(2 downto 0);
 signal SwRegister_sw_vcmd_axi_clk_gate_disable : std_logic;
 signal SwRegister_sw_vcmd_master_out_clk_gate_disable : std_logic;
 signal SwRegister_sw_vcmd_core_clk_gate_disable : std_logic;
 signal SwRegister_sw_vcmd_abort_mode : std_logic;
 signal SwRegister_sw_vcmd_reset_core : std_logic;
 signal SwRegister_sw_vcmd_reset_all : std_logic;
 signal SwRegister_sw_vcmd_start_trigger : std_logic;
 signal SwRegister_sw_vcmd_irq_intcmd : std_logic_vector(15 downto 0);
 signal SwRegister_sw_vcmd_irq_jmpp : std_logic;
 signal SwRegister_sw_vcmd_irq_jmpd : std_logic;
 signal SwRegister_sw_vcmd_irq_reset : std_logic;
 signal SwRegister_sw_vcmd_irq_abort : std_logic;
 signal SwRegister_sw_vcmd_irq_cmderr : std_logic;
 signal SwRegister_sw_vcmd_irq_timeout : std_logic;
 signal SwRegister_sw_vcmd_irq_buserr : std_logic;
 signal SwRegister_sw_vcmd_irq_endcmd : std_logic;
 signal SwRegister_sw_vcmd_irq_intcmd_en : std_logic_vector(15 downto 0);
 signal SwRegister_sw_vcmd_irq_jmpp_en : std_logic;
 signal SwRegister_sw_vcmd_irq_jmpd_en : std_logic;
 signal SwRegister_sw_vcmd_irq_reset_en : std_logic;
 signal SwRegister_sw_vcmd_irq_abort_en : std_logic;
 signal SwRegister_sw_vcmd_irq_cmderr_en : std_logic;
 signal SwRegister_sw_vcmd_irq_timeout_en : std_logic;
 signal SwRegister_sw_vcmd_irq_buserr_en : std_logic;
 signal SwRegister_sw_vcmd_irq_endcmd_en : std_logic;
 signal SwRegister_sw_vcmd_timeout_en : std_logic;
 signal SwRegister_sw_vcmd_timeout_cycles : std_logic_vector(30 downto 0);
 signal SwRegister_sw_vcmd_executing_cmd_addr : std_logic_vector(31 downto 0);
 signal SwRegister_sw_vcmd_executing_cmd_addr_msb : std_logic_vector(31 downto 0);
 signal SwRegister_sw_vcmd_exe_cmdbuf_length : std_logic_vector(15 downto 0);
 signal SwRegister_sw_vcmd_cmd_swap : std_logic_vector(3 downto 0);
 signal SwRegister_sw_vcmd_max_burst_len : std_logic_vector(7 downto 0);
 signal SwRegister_sw_vcmd_axi_id_rd : std_logic_vector(7 downto 0);
 signal SwRegister_sw_vcmd_axi_id_wr : std_logic_vector(7 downto 0);
 signal SwRegister_sw_vcmd_rdy_cmdbuf_count : std_logic_vector(31 downto 0);
 signal SwRegister_sw_vcmd_ext_abn_int_src_vcd_mmu_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_abn_int_src_vcd_l2cache_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_abn_int_src_vcd_dec400_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_abn_int_src_vcd_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_abn_int_src_cutree_mmu_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_abn_int_src_vce_mmu_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_abn_int_src_vce_l2cache_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_abn_int_src_vce_dec400_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_abn_int_src_cutree_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_abn_int_src_vce_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_vcd_mmu_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_vcd_l2cache_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_vcd_dec400_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_vcd_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_cutree_mmu_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_vce_mmu_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_vce_l2cache_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_vce_dec400_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_cutree_gate : std_logic;
 signal SwRegister_sw_vcmd_ext_norm_int_src_vce_gate : std_logic;
 signal SwRegister_sw_vcmd_cmdbuf_executing_id : std_logic_vector(31 downto 0);
