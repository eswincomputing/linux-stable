--register to signal map table from Document Version 1.1.2
 SwRegister_sw_vcmd_hw_id  <= swreg0(31 downto 16);
 SwRegister_sw_vcmd_hw_version  <= swreg0(15 downto 0);
 SwRegister_sw_vcmd_hw_build_date  <= swreg1(31 downto 0);
 SwRegister_sw_vcmd_ext_abn_int_src_vcd_mmu  <= swreg2(27);
 SwRegister_sw_vcmd_ext_abn_int_src_vcd_l2cache  <= swreg2(26);
 SwRegister_sw_vcmd_ext_abn_int_src_vcd_dec400  <= swreg2(25);
 SwRegister_sw_vcmd_ext_abn_int_src_vcd  <= swreg2(24);
 SwRegister_sw_vcmd_ext_abn_int_src_cutree_mmu  <= swreg2(21);
 SwRegister_sw_vcmd_ext_abn_int_src_vce_mmu  <= swreg2(20);
 SwRegister_sw_vcmd_ext_abn_int_src_vce_l2cache  <= swreg2(19);
 SwRegister_sw_vcmd_ext_abn_int_src_vce_dec400  <= swreg2(18);
 SwRegister_sw_vcmd_ext_abn_int_src_cutree  <= swreg2(17);
 SwRegister_sw_vcmd_ext_abn_int_src_vce  <= swreg2(16);
 SwRegister_sw_vcmd_ext_norm_int_src_vcd_mmu  <= swreg2(11);
 SwRegister_sw_vcmd_ext_norm_int_src_vcd_l2cache  <= swreg2(10);
 SwRegister_sw_vcmd_ext_norm_int_src_vcd_dec400  <= swreg2(9);
 SwRegister_sw_vcmd_ext_norm_int_src_vcd  <= swreg2(8);
 SwRegister_sw_vcmd_ext_norm_int_src_cutree_mmu  <= swreg2(5);
 SwRegister_sw_vcmd_ext_norm_int_src_vce_mmu  <= swreg2(4);
 SwRegister_sw_vcmd_ext_norm_int_src_vce_l2cache  <= swreg2(3);
 SwRegister_sw_vcmd_ext_norm_int_src_vce_dec400  <= swreg2(2);
 SwRegister_sw_vcmd_ext_norm_int_src_cutree  <= swreg2(1);
 SwRegister_sw_vcmd_ext_norm_int_src_vce  <= swreg2(0);
 SwRegister_sw_vcmd_exe_cmdbuf_count  <= swreg3(31 downto 0);
 SwRegister_sw_vcmd_executing_cmd  <= swreg4(31 downto 0);
 SwRegister_sw_vcmd_executing_cmd_msb  <= swreg5(31 downto 0);
 SwRegister_sw_vcmd_axi_total_ar_len  <= swreg6(31 downto 0);
 SwRegister_sw_vcmd_axi_total_r  <= swreg7(31 downto 0);
 SwRegister_sw_vcmd_axi_total_ar  <= swreg8(31 downto 0);
 SwRegister_sw_vcmd_axi_total_r_last  <= swreg9(31 downto 0);
 SwRegister_sw_vcmd_axi_total_aw_len  <= swreg10(31 downto 0);
 SwRegister_sw_vcmd_axi_total_w  <= swreg11(31 downto 0);
 SwRegister_sw_vcmd_axi_total_aw  <= swreg12(31 downto 0);
 SwRegister_sw_vcmd_axi_total_w_last  <= swreg13(31 downto 0);
 SwRegister_sw_vcmd_axi_total_b  <= swreg14(31 downto 0);
 SwRegister_sw_vcmd_axi_ar_valid  <= swreg15(31);
 SwRegister_sw_vcmd_axi_ar_ready  <= swreg15(30);
 SwRegister_sw_vcmd_axi_r_valid  <= swreg15(29);
 SwRegister_sw_vcmd_axi_r_ready  <= swreg15(28);
 SwRegister_sw_vcmd_axi_aw_valid  <= swreg15(27);
 SwRegister_sw_vcmd_axi_aw_ready  <= swreg15(26);
 SwRegister_sw_vcmd_axi_w_valid  <= swreg15(25);
 SwRegister_sw_vcmd_axi_w_ready  <= swreg15(24);
 SwRegister_sw_vcmd_axi_b_valid  <= swreg15(23);
 SwRegister_sw_vcmd_axi_b_ready  <= swreg15(22);
 SwRegister_sw_vcmd_work_state  <= swreg15(2 downto 0);
 SwRegister_sw_vcmd_axi_clk_gate_disable  <= swreg16(6);
 SwRegister_sw_vcmd_master_out_clk_gate_disable  <= swreg16(5);
 SwRegister_sw_vcmd_core_clk_gate_disable  <= swreg16(4);
 SwRegister_sw_vcmd_abort_mode  <= swreg16(3);
 SwRegister_sw_vcmd_reset_core  <= swreg16(2);
 SwRegister_sw_vcmd_reset_all  <= swreg16(1);
 SwRegister_sw_vcmd_start_trigger  <= swreg16(0);
 SwRegister_sw_vcmd_irq_intcmd  <= swreg17(31 downto 16);
 SwRegister_sw_vcmd_irq_jmpp  <= swreg17(7);
 SwRegister_sw_vcmd_irq_jmpd  <= swreg17(6);
 SwRegister_sw_vcmd_irq_reset  <= swreg17(5);
 SwRegister_sw_vcmd_irq_abort  <= swreg17(4);
 SwRegister_sw_vcmd_irq_cmderr  <= swreg17(3);
 SwRegister_sw_vcmd_irq_timeout  <= swreg17(2);
 SwRegister_sw_vcmd_irq_buserr  <= swreg17(1);
 SwRegister_sw_vcmd_irq_endcmd  <= swreg17(0);
 SwRegister_sw_vcmd_irq_intcmd_en  <= swreg18(31 downto 16);
 SwRegister_sw_vcmd_irq_jmpp_en  <= swreg18(7);
 SwRegister_sw_vcmd_irq_jmpd_en  <= swreg18(6);
 SwRegister_sw_vcmd_irq_reset_en  <= swreg18(5);
 SwRegister_sw_vcmd_irq_abort_en  <= swreg18(4);
 SwRegister_sw_vcmd_irq_cmderr_en  <= swreg18(3);
 SwRegister_sw_vcmd_irq_timeout_en  <= swreg18(2);
 SwRegister_sw_vcmd_irq_buserr_en  <= swreg18(1);
 SwRegister_sw_vcmd_irq_endcmd_en  <= swreg18(0);
 SwRegister_sw_vcmd_timeout_en  <= swreg19(31);
 SwRegister_sw_vcmd_timeout_cycles  <= swreg19(30 downto 0);
 SwRegister_sw_vcmd_executing_cmd_addr  <= swreg20(31 downto 0);
 SwRegister_sw_vcmd_executing_cmd_addr_msb  <= swreg21(31 downto 0);
 SwRegister_sw_vcmd_exe_cmdbuf_length  <= swreg22(15 downto 0);
 SwRegister_sw_vcmd_cmd_swap  <= swreg23(31 downto 28);
 SwRegister_sw_vcmd_max_burst_len  <= swreg23(23 downto 16);
 SwRegister_sw_vcmd_axi_id_rd  <= swreg23(15 downto 8);
 SwRegister_sw_vcmd_axi_id_wr  <= swreg23(7 downto 0);
 SwRegister_sw_vcmd_rdy_cmdbuf_count  <= swreg24(31 downto 0);
 SwRegister_sw_vcmd_ext_abn_int_src_vcd_mmu_gate  <= swreg25(28);
 SwRegister_sw_vcmd_ext_abn_int_src_vcd_l2cache_gate  <= swreg25(27);
 SwRegister_sw_vcmd_ext_abn_int_src_vcd_dec400_gate  <= swreg25(26);
 SwRegister_sw_vcmd_ext_abn_int_src_vcd_gate  <= swreg25(24);
 SwRegister_sw_vcmd_ext_abn_int_src_cutree_mmu_gate  <= swreg25(21);
 SwRegister_sw_vcmd_ext_abn_int_src_vce_mmu_gate  <= swreg25(20);
 SwRegister_sw_vcmd_ext_abn_int_src_vce_l2cache_gate  <= swreg25(19);
 SwRegister_sw_vcmd_ext_abn_int_src_vce_dec400_gate  <= swreg25(18);
 SwRegister_sw_vcmd_ext_abn_int_src_cutree_gate  <= swreg25(17);
 SwRegister_sw_vcmd_ext_abn_int_src_vce_gate  <= swreg25(16);
 SwRegister_sw_vcmd_ext_norm_int_src_vcd_mmu_gate  <= swreg25(11);
 SwRegister_sw_vcmd_ext_norm_int_src_vcd_l2cache_gate  <= swreg25(10);
 SwRegister_sw_vcmd_ext_norm_int_src_vcd_dec400_gate  <= swreg25(9);
 SwRegister_sw_vcmd_ext_norm_int_src_vcd_gate  <= swreg25(8);
 SwRegister_sw_vcmd_ext_norm_int_src_cutree_mmu_gate  <= swreg25(5);
 SwRegister_sw_vcmd_ext_norm_int_src_vce_mmu_gate  <= swreg25(4);
 SwRegister_sw_vcmd_ext_norm_int_src_vce_l2cache_gate  <= swreg25(3);
 SwRegister_sw_vcmd_ext_norm_int_src_vce_dec400_gate  <= swreg25(2);
 SwRegister_sw_vcmd_ext_norm_int_src_cutree_gate  <= swreg25(1);
 SwRegister_sw_vcmd_ext_norm_int_src_vce_gate  <= swreg25(0);
 SwRegister_sw_vcmd_cmdbuf_executing_id  <= swreg26(31 downto 0);
